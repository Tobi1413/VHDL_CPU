-------------------------------------------------------------------------------------------------------------
-- Project: VHDL_CPU
-- Author: Maher Popal & Tobias Blumers 
-- Description: 
-- Additional Comments:
-------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.riscv_types.all;

package program is
--  constant init_data_0 : ram_t := ("00000000", others => (others => '0'));
--  constant init_data_1 : ram_t := ("01010100", others => (others => '0'));
--  constant init_data_2 : ram_t := ("00000100", others => (others => '0'));
--  constant init_data_3 : ram_t := ("00010011", others => (others => '0'));
--  constant init_data_0 : ram_t := ("00000000", "00000000", "00000000", others => (others => '0'));
--  constant init_data_1 : ram_t := ("01010100", "01110100", "10010100", others => (others => '0'));
--  constant init_data_2 : ram_t := ("00000100", "10000100", "00000101", others => (others => '0'));
--  constant init_data_3 : ram_t := ("00010011", "10010011", "00110011", others => (others => '0'));
  
  

end program;

package body program is
end program;